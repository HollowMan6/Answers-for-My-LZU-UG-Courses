`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/05/24 16:31:55
// Design Name: 
// Module Name: BRAM_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SA4_CACHE_tb(

   );
reg clk;
reg rst;
reg[31:0] address;
   
SA4_CACHE SA4_CACHE_test(.clk(clk),.rst(rst),.address(address));

initial begin
rst = 1'b1;
clk = 1'b0;
address = 1'b0;
#5 rst = 1'b0;
#10 rst = 1'b1;
#5 clk =~clk;
   address <= 32'h1fffff50;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff58;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff88;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff90;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff98;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffa0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffa8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffb0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffb8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffc0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffc8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffd0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffd8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffe0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffffe8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1ffffff0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1ffffff8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000000;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000008;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000010;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000018;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000020;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000028;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000030;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000038;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000040;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000048;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000050;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000058;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000060;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000068;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000070;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000078;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000080;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000088;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000090;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h20000098;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000a0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000a8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000b0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000b8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000c0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000c8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000d0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000d8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000e0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000e8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000f0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h200000f8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h30031f10;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d960;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d968;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004caa0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d970;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d980;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h30000008;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d970;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d960;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d968;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004caa0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d978;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff58;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d978;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff68;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff68;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d980;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h30000008;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d970;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d960;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d968;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004caa0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d978;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff58;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d978;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff40;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff38;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff40;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff38;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff48;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h10034dc0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h0ffe7448;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h10034db0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h10034da0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h10034da8;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h10033ee0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d978;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff68;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004d978;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff78;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff78;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff78;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff78;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff30;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff28;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h3004cad0;
#5 clk =~clk;
#5 clk =~clk;
   address <= 32'h1fffff28;
#5 clk =~clk;
end

endmodule
